module uart (
    input i_Clk,
    input s_Tx,
    output u_Tx,
);
    reg u_Tx = 32'b0;
    reg u_Rx = 32'b0;
    
endmodule